
module compare(
			less,	//(input)
			equal,	//(input)
			comp 	//(output)
			);